// Code your testbench here
// or browse Examples
`include "tb_top.sv"
`include "test.sv"
